localparam [(NUM_COEFFS/2)*COEFF_WIDTH-1:0] COEFFS_VEC = 
1024'h0005_0007_000A_000E_0011_0016_001B_0021_0028_0030_0039_0044_0050_005E_006E_007F_0092_00A7_00BE_00D7_00F3_0110_0130_0152_0176_019C_01C4_01EF_021B_0249_0279_02AB_02DF_0313_0349_0381_03B9_03F2_042B_0465_049F_04D8_0512_054B_0583_05BA_05F0_0624_0657_0687_06B6_06E2_070C_0732_0756_0777_0795_07AF_07C6_07D9_07E8_07F4_07FC_07FF;