localparam [NUM_SLICES*COEFF_WIDTH-1:0] COEFFS_VEC = 
1024'h03FF_03FE_03FB_03F6_03F0_03E8_03DE_03D4_03C7_03BA_03AB_039A_0389_0376_0363_034E_0338_0322_030B_02F3_02DA_02C1_02A8_028E_0274_025A_023F_0225_020B_01F1_01D7_01BE_01A4_018C_0174_015C_0145_012F_011A_0105_00F1_00DE_00CC_00BB_00AB_009C_008D_0080_0074_0068_005E_0054_004B_0043_003C_0036_0030_002B_0027_0024_0021_001E_001D_001B;